/*~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
  SPI MODE 3
		CHANGE DATA @ NEGEDGE
		read data @posedge

 RSTB-active low asyn reset, CLK-clock, T_RB=0-rx  1-TX, mlb=0-LSB 1st 1-msb 1st
 START=1- starts data transmission cdiv 0=clk/4 1=/8   2=/16  3=/32
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~*/
module spi_master( rstb, clk, mlb, start, tdat, cdiv, din, ss, sck, dout, done, rdata );
input rstb,clk,mlb,start;
input [9:0] tdat;  //transmit data
input [1:0] cdiv;  //clock divider
input din;
output reg ss; 
output reg sck; 
output reg dout; 
output reg done;
output reg [9:0] rdata; //received data

parameter idle = 2'b00;
parameter send = 2'b10; 
parameter finish = 2'b11; 
reg [1:0] cur, nxt;
reg [9:0] treg, rreg;
reg [3:0] nbit;
reg [4:0] mid, cnt;
reg shift, clr;

//FSM i/o
always @(start or cur or nbit) begin
	nxt = cur;
	clr = 0;  
	shift = 0; //ss = 0;
	case ( cur )
		idle: begin
			if ( start == 1) begin 
				case ( cdiv )
					2'b00: mid = 2;
					2'b01: mid = 4;
					2'b10: mid = 8;
					2'b11: mid = 16;
 				endcase
				shift = 1;
				done = 1'b0;
				nxt = send;	 
			end
		end // idle		
		send: begin
			ss = 0;
			if ( nbit != 10 ) begin 
				shift = 1;
			end
			else begin
				rdata = rreg;
        done = 1'b1;
				nxt = finish;
			end
		end // send
		finish: begin
			shift = 0;
			ss = 1;
			clr = 1;
			nxt = idle;
		end
		default: nxt = finish;
  endcase
end // always

//state transistion
always@(negedge clk or negedge rstb) begin
	if( rstb == 0 ) 
		cur <= finish;
	else 
		cur <= nxt;
end

//setup falling edge (shift dout) sample rising edge (read din)
always@( negedge clk or posedge clr) begin
	if ( clr == 1 ) begin
    cnt = 0; 
    sck = 1;
  end
  else begin
		if ( shift == 1 ) begin
			cnt = cnt + 1; 
	  	if( cnt == mid ) begin
	  		sck = ~sck;
				cnt = 0;
			end //mid
		end //shift
	end //rst
end //always

//sample @ rising edge (read din)
always@( posedge sck or posedge clr ) begin // or negedge rstb
	if ( clr == 1 )  begin
		nbit = 0;
		rreg = 10'h3FF;
	end
	else begin 
	  if ( mlb == 0 ) begin //LSB first, din@msb -> right shift
		  rreg = { din, rreg[9:1] };
    end 
		else begin //MSB first, din@lsb -> left shift
		  rreg = { rreg[8:0], din };
    end
		nbit = nbit + 1;
	end //rst
end //always

always@(negedge sck or posedge clr) begin
	if ( clr == 1) begin
	  treg = 10'h3FF;
    dout = 1;  
	end  
	else begin
		if( nbit == 0 ) begin //load data into TREG
			treg = tdat;
      dout = mlb ? treg[9]:treg[0];
		end //nbit_if
		else begin
			if( mlb == 0 ) begin //LSB first, shift right
			  treg = { 1'b1, treg[9:1]};
        dout = treg[0];
      end
			else begin  //MSB first shift LEFT
		  	treg = { treg[8:0], 1'b1};
        dout = treg[9];
      end
		end
	end //rst
end //always

endmodule
